*IRF840 MCE 4-2-96
*500V  8A .85 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF840   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .402
RS  30  3  22.2M
RG  20  2  18.7
CGS  2  3  1.18N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.54N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=1.04MEG ETA=2M VTO=3 KP=4.33)
.MODEL DCGD D (CJO=1.54N VJ=.6 M=.68)
.MODEL DSUB D (IS=33.2N N=1.5 RS=.156 BV=500 CJO=817P VJ=.8 M=.42 TT=460N)
.MODEL DLIM D (IS=100U)
.ENDS IRF840


