*IRFIZ14G MCE  12/11/97
*Ref: International Rectifier Product Digest '94
*60V 8A .15ohm Power MOSFET pkg:TO-220 2,3,1
*SYM=POWMOSN
.SUBCKT IRFIZ14G 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  70.2M
RS  40  3  4.75M
RG  20  2  149
CGS  2  3  231P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  293P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=3.1 KP=3.44)
.MODEL DCGD D (CJO=293P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=33.2N N=1.5 RS=47.5M BV=60 CJO=447P VJ=0.8 M=0.42 TT=263N)
.MODEL DLIM D (IS=100U)
.ENDS 


