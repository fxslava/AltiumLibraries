*IRFZ44S MCE  12/4/97
*Ref: International Rectifier Product Digest '94
*60V 50A .024ohm Power MOSFET pkg:D2PAK 2,1,3
*SYM=POWMOSN
.SUBCKT IRFZ44S  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  10.4M
RS  40  3  1.6M
RG  20  2  3
CGS  2  3  1.44N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.83N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=3.1 KP=21.5)
.MODEL DCGD D (CJO=1.83N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=208N N=1.5 RS=7.6M BV=60 CJO=2.79N VJ=0.8 M=0.42 TT=456N)
.MODEL DLIM D (IS=100U)
.ENDS 


