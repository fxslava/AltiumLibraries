*IRLD014 MCE  12/11/97
*Ref: International Rectifier Product Digest '94
*60V 2A .706ohm Power MOSFET pkg:DIP4 1,4,3
*SYM=POWMOSN
.SUBCKT IRLD014  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.334
RS  40  3  18.6M
RG  20  2  885
CGS  2  3  49P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  62.2P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=3.1 KP=0.732)
.MODEL DCGD D (CJO=62.2P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=7.06N N=1.5 RS=0.224 BV=60 CJO=94.9P VJ=0.8 M=0.42 TT=165N)
.MODEL DLIM D (IS=100U)
.ENDS 


