*IRF820 MCE 4-2-96
*500V  2.5A 3 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF820   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  1.42
RS  30  3  76M
RG  20  2  60
CGS  2  3  323P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  475P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=1.04MEG ETA=2M VTO=3 KP=1.3)
.MODEL DCGD D (CJO=475P VJ=.6 M=.68)
.MODEL DSUB D (IS=10.3N N=1.5 RS=.34 BV=500 CJO=236P VJ=.8 M=.42 TT=260N)
.MODEL DLIM D (IS=100U)
.ENDS IRF820


