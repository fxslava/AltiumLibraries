*IRF9630S MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*200V 6A .185ohm Power MOSFET pkg:D2PAK 2,1,3
.SUBCKT IRF9630S 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  86.7M
RS  40  3  5.62M
RG  20  2  195
CGS  2  3  187P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  238P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=417K THETA=58.1M ETA=2M VTO=-3.1 KP=2)
.MODEL DCGD D (CJO=238P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=27N N=1.5 RS=69.2M BV=200 CJO=363P VJ=0.8 M=0.42 TT=247N)
.MODEL DLIM D (IS=100U)
.ENDS 


