*IRFZ14 MCE 4-9-96
*60V  10A .2 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFZ14   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  94M
RS  30  3  6M
RG  20  2  18.4
CGS  2  3  271P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  372P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=125K ETA=2M VTO=3 KP=1.29)
.MODEL DCGD D (CJO=372P VJ=.6 M=.68)
.MODEL DSUB D (IS=41.5N N=1.5 RS=85M BV=60 CJO=563P VJ=.8 M=.42 TT=70N)
.MODEL DLIM D (IS=100U)
.ENDS IRFZ14


