*IRF9Z24  MCE  4-2-96
*60V  11A  .28 ohms HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF9Z24  10 20 40 40
*     TERMINALS:  D  G  S
*  60 Volt  11 Amp  .28 ohm  P-Channel Power MOSFET  04-02-1996
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .132
RS  30  3  8M
RG  20  2  13.6
CGS  2  3  505P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  834P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 THETA=60M VMAX=125K ETA=2M VTO=-3 KP=.4)
.MODEL DCGD D (CJO=834P VJ=.6 M=.68)
.MODEL DSUB D (IS=45.6N N=1.5 RS=.504 BV=60 CJO=1.26N VJ=.8 M=.42 TT=100N)
.MODEL DLIM D (IS=100U)
.ENDS IRF9Z24

