*IRF830 MCE 4-2-96
*500V  4.5A 1.5 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF830   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .711
RS  30  3  38.5M
RG  20  2  33.3
CGS  2  3  542P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  873P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=1.04MEG ETA=2M VTO=3 KP=2)
.MODEL DCGD D (CJO=873P VJ=.6 M=.68)
.MODEL DSUB D (IS=18.6N N=1.5 RS=.188 BV=500 CJO=395P VJ=.8 M=.42 TT=320N)
.MODEL DLIM D (IS=100U)
.ENDS IRF830


