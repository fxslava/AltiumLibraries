*IRFIP140 MCE  12/11/97
*Ref: International Rectifier Product Digest '94
*100V 23A .0522ohm Power MOSFET pkg:TO-247 2,3,1
*SYM=POWMOSN
.SUBCKT IRFIP140 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  23.8M
RS  40  3  2.3M
RG  20  2  19.1
CGS  2  3  663P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  841P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=208K THETA=58.1M ETA=2M VTO=3.1 KP=8.29)
.MODEL DCGD D (CJO=841P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=95.5N N=1.5 RS=17.4M BV=100 CJO=1.28N VJ=0.8 M=0.42 TT=361N)
.MODEL DLIM D (IS=100U)
.ENDS 


