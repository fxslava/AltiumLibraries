*IRFZ24 MCE 4-9-96
*60V  17A .1 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFZ24   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  46.5M
RS  30  3  3.5M
RG  20  2  20
CGS  2  3  561P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.01N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=125K ETA=2M VTO=3 KP=4.08)
.MODEL DCGD D (CJO=1.01N VJ=.6 M=.68)
.MODEL DSUB D (IS=70.5N N=1.5 RS=44.1M BV=60 CJO=1.2N VJ=.8 M=.42 TT=88N)
.MODEL DLIM D (IS=100U)
.ENDS IRFZ24


