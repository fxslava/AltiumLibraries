*IRFIP350 MCE  12/11/97
*Ref: International Rectifier Product Digest '94
*400V 11A .109ohm Power MOSFET pkg:TO-247 2,3,1
*SYM=POWMOSN
.SUBCKT IRFIP350 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  50.8M
RS  40  3  3.73M
RG  20  2  94.5
CGS  2  3  317P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  402P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=833K THETA=58.1M ETA=2M VTO=3.1 KP=3.09)
.MODEL DCGD D (CJO=402P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=45.7N N=1.5 RS=50M BV=400 CJO=614P VJ=0.8 M=0.42 TT=289N)
.MODEL DLIM D (IS=100U)
.ENDS 

