*IRF7203 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*20V 4A .279ohm Power MOSFET pkg:SMD8A(A:8,1,2)(B:6,3,4)
.SUBCKT IRF7203  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.132
RS  40  3  7.98M
RG  20  2  320
CGS  2  3  124P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  157P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=41.7K THETA=58.1M ETA=2M VTO=-3.1 KP=3.36)
.MODEL DCGD D (CJO=157P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=17.8N N=1.5 RS=83.7M BV=20 CJO=240P VJ=0.8 M=0.42 TT=218N)
.MODEL DLIM D (IS=100U)
.ENDS 

