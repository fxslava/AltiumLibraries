*IRFZ34 MCE 4-9-96
*60V  30A .05 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFZ34   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  22.7M
RS  30  3  2.25M
RG  20  2  19.4
CGS  2  3  1.1N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.28N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=125K ETA=2M VTO=3 KP=6.48)
.MODEL DCGD D (CJO=1.28N VJ=.6 M=.68)
.MODEL DSUB D (IS=124N N=1.5 RS=28.3M BV=60 CJO=2.15N VJ=.8 M=.42 TT=120N)
.MODEL DLIM D (IS=100U)
.ENDS IRFZ34


