*IRF9540  MCE  4-2-96
*100V  19A  .2 ohms HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF9540  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  94M
RS  30  3  6M
RG  20  2  17.6
CGS  2  3  1.26N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  1.79N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 THETA=60M VMAX=208K ETA=2M VTO=-3 KP=3.95)
.MODEL DCGD D (CJO=1.79N VJ=.6 M=.68)
.MODEL DSUB D (IS=78.9N N=1.5 RS=.223 BV=100 CJO=1.93N VJ=.8 M=.42 TT=130N)
.MODEL DLIM D (IS=100U)
.ENDS IRF9540


