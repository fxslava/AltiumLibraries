*IRFZ24S MCE  12/4/97
*Ref: International Rectifier Product Digest '94
*60V 17A .0706ohm Power MOSFET pkg:D2PAK 2,1,3
*SYM=POWMOSN
.SUBCKT IRFZ24S  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  32.5M
RS  40  3  2.76M
RG  20  2  43.5
CGS  2  3  490P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  622P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=3.1 KP=7.32)
.MODEL DCGD D (CJO=622P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=70.6N N=1.5 RS=22.4M BV=60 CJO=949P VJ=0.8 M=0.42 TT=330N)
.MODEL DLIM D (IS=100U)
.ENDS 


