*IRF9Z14S MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*60V 7A .179ohm Power MOSFET pkg:D2PAK 2,1,3
.SUBCKT IRF9Z14S 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  84.1M
RS  40  3  5.48M
RG  20  2  187
CGS  2  3  193P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  245P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=-3.1 KP=2.88)
.MODEL DCGD D (CJO=245P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=27.8N N=1.5 RS=56.7M BV=60 CJO=374P VJ=0.8 M=0.42 TT=249N)
.MODEL DLIM D (IS=100U)
.ENDS 


