*IRFIP9240 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*200V 9A .135ohm Power MOSFET pkg:TO-247 2,3,1
.SUBCKT IRFIP9240 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  63M
RS  40  3  4.37M
RG  20  2  129
CGS  2  3  256P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  326P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=417K THETA=58.1M ETA=2M VTO=-3.1 KP=2.74)
.MODEL DCGD D (CJO=326P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=36.9N N=1.5 RS=50.6M BV=200 CJO=497P VJ=0.8 M=0.42 TT=272N)
.MODEL DLIM D (IS=100U)
.ENDS 


