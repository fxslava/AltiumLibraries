*IRFL9014 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*60V 2A .667ohm Power MOSFET pkg:SOT-223 2,1,3
.SUBCKT IRFL9014 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.316
RS  40  3  17.7M
RG  20  2  833
CGS  2  3  51.9P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  65.9P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=-3.1 KP=0.775)
.MODEL DCGD D (CJO=65.9P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=7.47N N=1.5 RS=0.211 BV=60 CJO=101P VJ=0.8 M=0.42 TT=168N)
.MODEL DLIM D (IS=100U)
.ENDS 


