*IRFPG50 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*1000V 6A .197ohm Power MOSFET pkg:TO-247 2,3,1
*SYM=POWMOSN
.SUBCKT IRFPG50  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  92.4M
RS  40  3  5.92M
RG  20  2  211
CGS  2  3  176P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  223P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=1 LAMBDA=2M VTO=3.1 KP=1.37)
.MODEL DCGD D (CJO=223P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=25.3N N=1.5 RS=0.139 BV=1K CJO=341P VJ=0.8 M=0.42 TT=243N)
.MODEL DLIM D (IS=100U)
.ENDS 


