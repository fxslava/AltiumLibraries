*IRFPG42 MCE 5/21/98
*1000V  4A 4.2 ohm Power MOSFET pkg:TO-247 2,1,3
.SUBCKT IRFPG42  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  1.99
RS  40  3  0.106
RG  20  2  223
CGS  2  3  116P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  147P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=1 LAMBDA=2M VTO=3 KP=3.43)
.MODEL DCGD D (CJO=147P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=16.2N N=1.5 RS=0.269 BV=1K CJO=225P VJ=0.8 M=0.42 TT=1U)
.MODEL DLIM D (IS=100U)
.ENDS 


