*IRF9630  MCE  4-2-96
*200V  6.5A  .8 ohms HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF9630  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .379
RS  30  3  21M
RG  20  2  23
CGS  2  3  660P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  513P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 THETA=60M VMAX=416K ETA=2M VTO=-3 KP=1.94)
.MODEL DCGD D (CJO=513P VJ=.6 M=.68)
.MODEL DSUB D (IS=26.9N N=1.5 RS=.885 BV=200 CJO=688P VJ=.8 M=.42 TT=200N)
.MODEL DLIM D (IS=100U)
.ENDS IRF9630


