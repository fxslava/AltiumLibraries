*IRF734 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*450V 5A .245ohm Power MOSFET pkg:TO-220 2,3,1
*SYM=POWMOSN
.SUBCKT IRF734   10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.115
RS  40  3  7.12M
RG  20  2  274
CGS  2  3  141P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  179P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=937K THETA=58.1M ETA=2M VTO=3.1 KP=1.36)
.MODEL DCGD D (CJO=179P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=20.3N N=1.5 RS=0.117 BV=450 CJO=274P VJ=0.8 M=0.42 TT=227N)
.MODEL DLIM D (IS=100U)
.ENDS 

