*IRFS1Z0  MCE  12/2/97
*Ref: International Rectifier Product Digest '94
*100V 1A 1.46ohm Power MOSFET pkg:SOT-89 2,1,3
*SYM=POWMOSN
.SUBCKT IRFS1Z0  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.694
RS  40  3  37.6M
RG  20  2  1.89K
CGS  2  3  23.6P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  30P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=208K THETA=58.1M ETA=2M VTO=3.1 KP=0.295)
.MODEL DCGD D (CJO=30P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=3.4N N=1.5 RS=0.488 BV=100 CJO=45.8P VJ=0.8 M=0.42 TT=133N)
.MODEL DLIM D (IS=100U)
.ENDS 


