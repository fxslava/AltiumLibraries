*50V 15A .1 ohm  HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFZ20 10 20 30 30
M1   4  1  5  5  DMOS L=1U W=1U
RG  20  1  10
RD  10  4  37M
RDS  4  5  1.18MEG
CGD  7  4  590P
RCG  7  4  10MEG
MCG  7  9  1  1  SW
ECG  9  1  1  4  1
DGD  1  6  DCGD
MDG  6  8  4  4  SW
EDG  8  4  4  1  1
DDS  5  4  DSUB
LS   5 30  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=1.6MEG THETA=300M VTO=3.2
+ KP=5.0 RS=5M IS=2.16P CGSO=725U)
.MODEL SW   NMOS (LEVEL=3 VTO=0 KP=20)
.MODEL DCGD D (CJO=590P M=.5 VJ=.41)
.MODEL DSUB D (IS=2.16P RS=0 BV=50 IBV=.001
+ VJ=.8 M=.4 CJO=902P TT=144N)
.ENDS IRFZ20


