*IRF614 MCE 4-2-96
*250V  2.7A 2 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF614   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .949
RS  30  3  51M
RG  20  2  55.5
CGS  2  3  130P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  123P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=521K ETA=2M VTO=3 KP=.472)
.MODEL DCGD D (CJO=123P VJ=.6 M=.68)
.MODEL DSUB D (IS=11.2N N=1.5 RS=.463 BV=250 CJO=139P VJ=.8 M=.42 TT=190N)
.MODEL DLIM D (IS=100U)
.ENDS IRF614


