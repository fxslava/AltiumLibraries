*IRFK6JC50 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*600V 48A .025ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
.SUBCKT IRFK6JC50 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  10.9M
RS  40  3  1.62M
RG  20  2  3.12
CGS  2  3  1.38N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.76N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=1 LAMBDA=2M VTO=3.1 KP=10.8)
.MODEL DCGD D (CJO=1.76N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=199N N=1.5 RS=13.5M BV=600 IBV=5M CJO=2.68N VJ=0.8 M=0.42 TT=450N)
.MODEL DLIM D (IS=100U)
.ENDS 


