*IRF624 MCE 4-2-96
*250V  4.4A 1.1 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF624   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .521
RS  30  3  28.5M
RG  20  2  34.1
CGS  2  3  245P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  192P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=521K ETA=2M VTO=3 KP=.807)
.MODEL DCGD D (CJO=192P VJ=.6 M=.68)
.MODEL DSUB D (IS=18.2N N=1.5 RS=.238 BV=250 CJO=266P VJ=.8 M=.42 TT=200N)
.MODEL DLIM D (IS=100U)
.ENDS IRF624


