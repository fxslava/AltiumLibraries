*IRLR120 MCE  12/4/97
*Ref: International Rectifier Product Digest '94
*100V 8A .156ohm Power MOSFET pkg:DPAK 2,1,3
*SYM=POWMOSN
.SUBCKT IRLR120  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  73M
RS  40  3  4.9M
RG  20  2  156
CGS  2  3  222P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  282P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=208K THETA=58.1M ETA=2M VTO=3.1 KP=2.77)
.MODEL DCGD D (CJO=282P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=32N N=1.5 RS=51.9M BV=100 CJO=430P VJ=0.8 M=0.42 TT=260N)
.MODEL DLIM D (IS=100U)
.ENDS 


