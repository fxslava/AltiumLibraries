*IRFK4JC50 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*600V 35A .0343ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
.SUBCKT IRFK4JC50 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  15.3M
RS  40  3  1.86M
RG  20  2  4.29
CGS  2  3  1.01N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.28N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=1 LAMBDA=2M VTO=3.1 KP=7.84)
.MODEL DCGD D (CJO=1.28N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=145N N=1.5 RS=18.6M BV=600 IBV=4M CJO=1.95N VJ=0.8 M=0.42 TT=410N)
.MODEL DLIM D (IS=100U)
.ENDS 


