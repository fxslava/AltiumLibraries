*IRF9Z14  MCE  4-2-96
*60V  6.7A  .5 ohms HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF9Z14  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .236
RS  30  3  13.5M
RG  20  2  45.6
CGS  2  3  239P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  398P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 THETA=60M VMAX=125K ETA=2M VTO=-3 KP=.661)
.MODEL DCGD D (CJO=398P VJ=.6 M=.68)
.MODEL DSUB D (IS=27.8N N=1.5 RS=.709 BV=60 CJO=598P VJ=.8 M=.42 TT=80N)
.MODEL DLIM D (IS=100U)
.ENDS IRF9Z14


