*IRF710S MCE  12/4/97
*Ref: International Rectifier Product Digest '94
*400V 2A .6ohm Power MOSFET pkg:D2PAK 2,1,3
*SYM=POWMOSN
.SUBCKT IRF710S  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.284
RS  40  3  16M
RG  20  2  745
CGS  2  3  57.6P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  73.2P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=833K THETA=58.1M ETA=2M VTO=3.1 KP=0.563)
.MODEL DCGD D (CJO=73.2P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=8.3N N=1.5 RS=0.275 BV=400 CJO=112P VJ=0.8 M=0.42 TT=174N)
.MODEL DLIM D (IS=100U)
.ENDS 


