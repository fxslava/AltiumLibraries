* jjt 5/6/2000: deleted redundant first model 
* jjt 5/4/2002: changed sign of VTO to match PD-9.519E (CAPS) datasheet.
*IRFU9110 MCE  5/27/98
*100V 3A 1.2ohm Power MOSFET pkg:TO251AA 2,1,3
.SUBCKT IRFU9110 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.569
RS  40  3  31M
RG  20  2  48.4
CGS  2  3  272P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  231P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=208K THETA=60M ETA=2M VTO=-3 KP=1.2)
.MODEL DCGD D (CJO=231P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=12.9N N=1.5 RS=1.53 BV=100 CJO=327P VJ=0.8 M=0.42 TT=105N)
.MODEL DLIM D (IS=100U)
.ENDS 

* Origin: Mcemos.lib
