*IRFI9Z14G MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*60V 5A .226ohm Power MOSFET pkg:TO-220 2,3,1
.SUBCKT IRFI9Z14G 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.107
RS  40  3  6.66M
RG  20  2  250
CGS  2  3  153P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  194P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=-3.1 KP=2.28)
.MODEL DCGD D (CJO=194P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=22N N=1.5 RS=71.7M BV=60 CJO=296P VJ=0.8 M=0.42 TT=233N)
.MODEL DLIM D (IS=100U)
.ENDS 


