*IRF740 MCE 4-2-96
*400V  10A .55 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF740   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .26
RS  30  3  14.7M
RG  20  2  15
CGS  2  3  1.28N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.54N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=833K ETA=2M VTO=3 KP=4.95)
.MODEL DCGD D (CJO=1.54N VJ=.6 M=.68)
.MODEL DSUB D (IS=41.5N N=1.5 RS=.125 BV=400 CJO=903P VJ=.8 M=.42 TT=370N)
.MODEL DLIM D (IS=100U)
.ENDS IRF740


