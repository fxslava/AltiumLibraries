*IRFZ46 MCE 4-9-96
*50V  50A .024 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFZ46   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  10.4M
RS  30  3  1.6M
RG  20  2  27.8
CGS  2  3  1.64N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  2.05N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=104K ETA=2M VTO=3 KP=33.2)
.MODEL DCGD D (CJO=2.05N VJ=.6 M=.68)
.MODEL DSUB D (IS=207N N=1.5 RS=35M BV=50 CJO=3.44N VJ=.8 M=.42 TT=66N)
.MODEL DLIM D (IS=100U)
.ENDS IRFZ46


