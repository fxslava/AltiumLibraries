*IRF710 MCE 4-2-96
*400V  2A 3.6 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF710   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  1.7
RS  30  3  91M
RG  20  2  75
CGS  2  3  163P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  80.9P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=833K ETA=2M VTO=3 KP=.736)
.MODEL DCGD D (CJO=80.9P VJ=.6 M=.68)
.MODEL DSUB D (IS=8.3N N=1.5 RS=.425 BV=400 CJO=119P VJ=.8 M=.42 TT=240N)
.MODEL DLIM D (IS=100U)
.ENDS IRF710


