*IRFBF20 MCE 4-9-96
*900V 1.7A 8 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFBF20  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  3.8
RS  30  3  .201
RG  20  2  88.2
CGS  2  3  472P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  231P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=1 LAMBDA=2M VTO=3 KP=.252)
.MODEL DCGD D (CJO=231P VJ=.6 M=.68)
.MODEL DSUB D (IS=7.05N N=1.5 RS=.441 BV=900 CJO=159P VJ=.8 M=.42 TT=350N)
.MODEL DLIM D (IS=100U)
.ENDS IRFBF20


