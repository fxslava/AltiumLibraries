*IRF9530
*Harris P-ch. BVdss=100V Ids=12A Rds(on)=.3 ohms: D G S
.SUBCKT IRF9530 10 20 30 30
M1   4  1  5  5  DMOS L=1U W=1U
RG  20  1  21.4
RD  10  4  .117
RDS  4  5  2.54MEG
CGD  7  4  787P
RCG  7  4  10MEG
MCG  7  9  1  1  SW
ECG  9  1  1  4  1
DGD  6  1  DCGD
MDG  6  8  4  4  SW
EDG  8  4  4  1  1
DDS  4  5  DSUB
LS   5 30  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=6.6MEG THETA=220M VTO=-3.2
+ KP=3.2 RS=8.25M IS=504F CGSO=400U)
.MODEL SW   PMOS (LEVEL=3 VTO=0 KP=20)
.MODEL DCGD D (CJO=787P M=.5 VJ=.41)
.MODEL DSUB D (IS=504F RS=.513 BV=100 IBV=.001
+ VJ=.8 M=.4 CJO=802P TT=432N)
.ENDS IRF9530


