*IRFZ48 MCE 4-8-96
*60V  50A .018 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRFZ48   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  7.55M
RS  30  3  1.45M
RG  20  2  68.4
CGS  2  3  2.21N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  2.44N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=125K ETA=2M VTO=3 KP=22.8)
.MODEL DCGD D (CJO=2.44N VJ=.6 M=.68)
.MODEL DSUB D (IS=207N N=1.5 RS=25M BV=60 CJO=4.77N VJ=.8 M=.42 TT=120N)
.MODEL DLIM D (IS=100U)
.ENDS IRFZ48


