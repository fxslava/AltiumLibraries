*IRF7102 MCE 4-2-96
*50V  2A .3 ohm HEXFET pkg:SO-8 (A:8,2,1)(B:6,4,3)
.SUBCKT IRF7102  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .141
RS  30  3  8.5M
RG  20  2  75
CGS  2  3  108P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  154P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  6N
.MODEL DMOS NMOS (LEVEL=3 THETA=80M VMAX=104K ETA=2M VTO=2.25 KP=1)
.MODEL DCGD D (CJO=154P VJ=.6 M=.68)
.MODEL DSUB D (IS=8.3N N=1.5 RS=.325 BV=50 CJO=219P VJ=.8 M=.42 TT=38N)
.MODEL DLIM D (IS=100U)
.ENDS IRF7102


