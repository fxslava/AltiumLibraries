* jjt 5/6/2000: deleted redundant first model 

*IRFU9220 MCE  5/27/98
*200V 4A 1.5ohm Power MOSFET pkg:TO251AA 2,1,3
.SUBCKT IRFU9220 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.712
RS  40  3  38.5M
RG  20  2  41.7
CGS  2  3  517P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  424P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=417K THETA=60M ETA=2M VTO=-3 KP=1.19)
.MODEL DCGD D (CJO=424P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=14.9N N=1.5 RS=1.54 BV=200 CJO=331P VJ=0.8 M=0.42 TT=150N)
.MODEL DLIM D (IS=100U)
.ENDS 

* Origin: Mcemos.lib
