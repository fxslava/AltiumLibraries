*IRF644 MCE 4-2-96
*250V  14A .28 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF644   10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .132
RS  30  3  8M
RG  20  2  21.6
CGS  2  3  1.21N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.09N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=521K ETA=2M VTO=3 KP=4.98)
.MODEL DCGD D (CJO=1.09N VJ=.6 M=.68)
.MODEL DSUB D (IS=58.1N N=1.5 RS=75M BV=250 CJO=1.05N VJ=.8 M=.42 TT=250N)
.MODEL DLIM D (IS=100U)
.ENDS IRF644


