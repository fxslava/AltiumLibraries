*IRFK6J350 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*400V 75A .016ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
.SUBCKT IRFK6J350 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  6.6M
RS  40  3  1.4M
RG  20  2  2
CGS  2  3  2.16N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  2.74N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=833K THETA=58.1M ETA=2M VTO=3.1 KP=21.1)
.MODEL DCGD D (CJO=2.74N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=311N N=1.5 RS=7.33M BV=400 IBV=5M CJO=4.19N VJ=0.8 M=0.42 TT=515N)
.MODEL DLIM D (IS=100U)
.ENDS 


