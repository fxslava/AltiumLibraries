*IRF530 MCE 2-20-96
*100V  14A .16 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF530  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  39.7M
RS  30  3  3.14M
RG  20  2  13
CGS  2  3  610P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  770P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=208K ETA=2M VTO=3 KP=4.5)
.MODEL DCGD D (CJO=770P VJ=.6 M=.68)
.MODEL DSUB D (IS=58.1N N=1.5 RS=28.5M BV=100 CJO=817P VJ=.8 M=.42 TT=150N)
.MODEL DLIM D (IS=100U)
.ENDS IRF530


