*IRLS0Z0  MCE  12/2/97
*Ref: International Rectifier Product Digest '94
*50V 3A .462ohm Power MOSFET pkg:SOT-89 2,1,3
*SYM=POWMOSN
.SUBCKT IRLS0Z0  10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.218
RS  40  3  12.5M
RG  20  2  561
CGS  2  3  74.9P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  95.1P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=104K THETA=58.1M ETA=2M VTO=3.1 KP=1.21)
.MODEL DCGD D (CJO=95.1P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=10.8N N=1.5 RS=0.144 BV=50 CJO=145P VJ=0.8 M=0.42 TT=188N)
.MODEL DLIM D (IS=100U)
.ENDS 


