* jjt 5/6/2000: deleted redundant first model 

*IRFU9120 MCE  5/27/98
*100V 6A .6ohm Power MOSFET pkg:TO251AA 2,1,3
.SUBCKT IRFU9120 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  0.284
RS  40  3  16M
RG  20  2  26.8
CGS  2  3  440P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  578P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=208K THETA=60M ETA=2M VTO=-3 KP=2.16)
.MODEL DCGD D (CJO=578P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=23.2N N=1.5 RS=0.991 BV=100 CJO=538P VJ=0.8 M=0.42 TT=130N)
.MODEL DLIM D (IS=100U)
.ENDS 

* Origin: Mcemos.lib