*IRF9620  MCE  4-2-96
*200V  3.5A  1.5 ohms HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF9620  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .711
RS  30  3  38.5M
RG  20  2  42.8
CGS  2  3  320P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  385P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 THETA=60M VMAX=416K ETA=2M VTO=-3 KP=.643)
.MODEL DCGD D (CJO=385P VJ=.6 M=.68)
.MODEL DSUB D (IS=14.5N N=1.5 RS=1.78 BV=200 CJO=301P VJ=.8 M=.42 TT=300N)
.MODEL DLIM D (IS=100U)
.ENDS IRF9620


